// QsysSystem.v

// Generated using ACDS version 16.1 196

`timescale 1 ps / 1 ps
module QsysSystem (
		input  wire        clk_clk,                                    //                                 clk.clk
		output wire [7:0]  green_leds_external_connection_export,      //      green_leds_external_connection.export
		input  wire [3:0]  keys_external_connection_export,            //            keys_external_connection.export
		output wire [17:0] red_leds_external_connection_export,        //        red_leds_external_connection.export
		input  wire        reset_reset,                                //                               reset.reset
		output wire        sdram_clk_clk,                              //                           sdram_clk.clk
		output wire [12:0] sdram_wire_addr,                            //                          sdram_wire.addr
		output wire [1:0]  sdram_wire_ba,                              //                                    .ba
		output wire        sdram_wire_cas_n,                           //                                    .cas_n
		output wire        sdram_wire_cke,                             //                                    .cke
		output wire        sdram_wire_cs_n,                            //                                    .cs_n
		inout  wire [31:0] sdram_wire_dq,                              //                                    .dq
		output wire [3:0]  sdram_wire_dqm,                             //                                    .dqm
		output wire        sdram_wire_ras_n,                           //                                    .ras_n
		output wire        sdram_wire_we_n,                            //                                    .we_n
		output wire [31:0] sevseg4msb_external_connection_export,      //      sevseg4msb_external_connection.export
		output wire [31:0] sevsegment_4lsb_external_connection_export, // sevsegment_4lsb_external_connection.export
		input  wire [17:0] switches_external_connection_export         //        switches_external_connection.export
	);

	wire         clk_sys_clk_clk;                                           // CLK:sys_clk_clk -> [GREEN_LEDs:clk, JTAG_UART:clk, KEYS:clk, On_Chip_Mem:clk, Processor:clk, RED_LEDs:clk, SDRAM:clk, SYSID:clock, SevSeg4MSB:clk, SevSegment_4LSB:clk, Switches:clk, irq_mapper:clk, mm_interconnect_0:CLK_sys_clk_clk, rst_controller:clk, timer_0:clk, timer_1:clk]
	wire  [31:0] processor_data_master_readdata;                            // mm_interconnect_0:Processor_data_master_readdata -> Processor:d_readdata
	wire         processor_data_master_waitrequest;                         // mm_interconnect_0:Processor_data_master_waitrequest -> Processor:d_waitrequest
	wire         processor_data_master_debugaccess;                         // Processor:jtag_debug_module_debugaccess_to_roms -> mm_interconnect_0:Processor_data_master_debugaccess
	wire  [28:0] processor_data_master_address;                             // Processor:d_address -> mm_interconnect_0:Processor_data_master_address
	wire   [3:0] processor_data_master_byteenable;                          // Processor:d_byteenable -> mm_interconnect_0:Processor_data_master_byteenable
	wire         processor_data_master_read;                                // Processor:d_read -> mm_interconnect_0:Processor_data_master_read
	wire         processor_data_master_readdatavalid;                       // mm_interconnect_0:Processor_data_master_readdatavalid -> Processor:d_readdatavalid
	wire         processor_data_master_write;                               // Processor:d_write -> mm_interconnect_0:Processor_data_master_write
	wire  [31:0] processor_data_master_writedata;                           // Processor:d_writedata -> mm_interconnect_0:Processor_data_master_writedata
	wire  [31:0] processor_instruction_master_readdata;                     // mm_interconnect_0:Processor_instruction_master_readdata -> Processor:i_readdata
	wire         processor_instruction_master_waitrequest;                  // mm_interconnect_0:Processor_instruction_master_waitrequest -> Processor:i_waitrequest
	wire  [28:0] processor_instruction_master_address;                      // Processor:i_address -> mm_interconnect_0:Processor_instruction_master_address
	wire         processor_instruction_master_read;                         // Processor:i_read -> mm_interconnect_0:Processor_instruction_master_read
	wire         processor_instruction_master_readdatavalid;                // mm_interconnect_0:Processor_instruction_master_readdatavalid -> Processor:i_readdatavalid
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect;  // mm_interconnect_0:JTAG_UART_avalon_jtag_slave_chipselect -> JTAG_UART:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata;    // JTAG_UART:av_readdata -> mm_interconnect_0:JTAG_UART_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest; // JTAG_UART:av_waitrequest -> mm_interconnect_0:JTAG_UART_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_address;     // mm_interconnect_0:JTAG_UART_avalon_jtag_slave_address -> JTAG_UART:av_address
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;        // mm_interconnect_0:JTAG_UART_avalon_jtag_slave_read -> JTAG_UART:av_read_n
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;       // mm_interconnect_0:JTAG_UART_avalon_jtag_slave_write -> JTAG_UART:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata;   // mm_interconnect_0:JTAG_UART_avalon_jtag_slave_writedata -> JTAG_UART:av_writedata
	wire  [31:0] mm_interconnect_0_sysid_control_slave_readdata;            // SYSID:readdata -> mm_interconnect_0:SYSID_control_slave_readdata
	wire   [0:0] mm_interconnect_0_sysid_control_slave_address;             // mm_interconnect_0:SYSID_control_slave_address -> SYSID:address
	wire  [31:0] mm_interconnect_0_processor_jtag_debug_module_readdata;    // Processor:jtag_debug_module_readdata -> mm_interconnect_0:Processor_jtag_debug_module_readdata
	wire         mm_interconnect_0_processor_jtag_debug_module_waitrequest; // Processor:jtag_debug_module_waitrequest -> mm_interconnect_0:Processor_jtag_debug_module_waitrequest
	wire         mm_interconnect_0_processor_jtag_debug_module_debugaccess; // mm_interconnect_0:Processor_jtag_debug_module_debugaccess -> Processor:jtag_debug_module_debugaccess
	wire   [8:0] mm_interconnect_0_processor_jtag_debug_module_address;     // mm_interconnect_0:Processor_jtag_debug_module_address -> Processor:jtag_debug_module_address
	wire         mm_interconnect_0_processor_jtag_debug_module_read;        // mm_interconnect_0:Processor_jtag_debug_module_read -> Processor:jtag_debug_module_read
	wire   [3:0] mm_interconnect_0_processor_jtag_debug_module_byteenable;  // mm_interconnect_0:Processor_jtag_debug_module_byteenable -> Processor:jtag_debug_module_byteenable
	wire         mm_interconnect_0_processor_jtag_debug_module_write;       // mm_interconnect_0:Processor_jtag_debug_module_write -> Processor:jtag_debug_module_write
	wire  [31:0] mm_interconnect_0_processor_jtag_debug_module_writedata;   // mm_interconnect_0:Processor_jtag_debug_module_writedata -> Processor:jtag_debug_module_writedata
	wire         mm_interconnect_0_on_chip_mem_s1_chipselect;               // mm_interconnect_0:On_Chip_Mem_s1_chipselect -> On_Chip_Mem:chipselect
	wire  [31:0] mm_interconnect_0_on_chip_mem_s1_readdata;                 // On_Chip_Mem:readdata -> mm_interconnect_0:On_Chip_Mem_s1_readdata
	wire   [9:0] mm_interconnect_0_on_chip_mem_s1_address;                  // mm_interconnect_0:On_Chip_Mem_s1_address -> On_Chip_Mem:address
	wire   [3:0] mm_interconnect_0_on_chip_mem_s1_byteenable;               // mm_interconnect_0:On_Chip_Mem_s1_byteenable -> On_Chip_Mem:byteenable
	wire         mm_interconnect_0_on_chip_mem_s1_write;                    // mm_interconnect_0:On_Chip_Mem_s1_write -> On_Chip_Mem:write
	wire  [31:0] mm_interconnect_0_on_chip_mem_s1_writedata;                // mm_interconnect_0:On_Chip_Mem_s1_writedata -> On_Chip_Mem:writedata
	wire         mm_interconnect_0_on_chip_mem_s1_clken;                    // mm_interconnect_0:On_Chip_Mem_s1_clken -> On_Chip_Mem:clken
	wire         mm_interconnect_0_red_leds_s1_chipselect;                  // mm_interconnect_0:RED_LEDs_s1_chipselect -> RED_LEDs:chipselect
	wire  [31:0] mm_interconnect_0_red_leds_s1_readdata;                    // RED_LEDs:readdata -> mm_interconnect_0:RED_LEDs_s1_readdata
	wire   [1:0] mm_interconnect_0_red_leds_s1_address;                     // mm_interconnect_0:RED_LEDs_s1_address -> RED_LEDs:address
	wire         mm_interconnect_0_red_leds_s1_write;                       // mm_interconnect_0:RED_LEDs_s1_write -> RED_LEDs:write_n
	wire  [31:0] mm_interconnect_0_red_leds_s1_writedata;                   // mm_interconnect_0:RED_LEDs_s1_writedata -> RED_LEDs:writedata
	wire         mm_interconnect_0_green_leds_s1_chipselect;                // mm_interconnect_0:GREEN_LEDs_s1_chipselect -> GREEN_LEDs:chipselect
	wire  [31:0] mm_interconnect_0_green_leds_s1_readdata;                  // GREEN_LEDs:readdata -> mm_interconnect_0:GREEN_LEDs_s1_readdata
	wire   [1:0] mm_interconnect_0_green_leds_s1_address;                   // mm_interconnect_0:GREEN_LEDs_s1_address -> GREEN_LEDs:address
	wire         mm_interconnect_0_green_leds_s1_write;                     // mm_interconnect_0:GREEN_LEDs_s1_write -> GREEN_LEDs:write_n
	wire  [31:0] mm_interconnect_0_green_leds_s1_writedata;                 // mm_interconnect_0:GREEN_LEDs_s1_writedata -> GREEN_LEDs:writedata
	wire         mm_interconnect_0_sevsegment_4lsb_s1_chipselect;           // mm_interconnect_0:SevSegment_4LSB_s1_chipselect -> SevSegment_4LSB:chipselect
	wire  [31:0] mm_interconnect_0_sevsegment_4lsb_s1_readdata;             // SevSegment_4LSB:readdata -> mm_interconnect_0:SevSegment_4LSB_s1_readdata
	wire   [1:0] mm_interconnect_0_sevsegment_4lsb_s1_address;              // mm_interconnect_0:SevSegment_4LSB_s1_address -> SevSegment_4LSB:address
	wire         mm_interconnect_0_sevsegment_4lsb_s1_write;                // mm_interconnect_0:SevSegment_4LSB_s1_write -> SevSegment_4LSB:write_n
	wire  [31:0] mm_interconnect_0_sevsegment_4lsb_s1_writedata;            // mm_interconnect_0:SevSegment_4LSB_s1_writedata -> SevSegment_4LSB:writedata
	wire  [31:0] mm_interconnect_0_switches_s1_readdata;                    // Switches:readdata -> mm_interconnect_0:Switches_s1_readdata
	wire   [1:0] mm_interconnect_0_switches_s1_address;                     // mm_interconnect_0:Switches_s1_address -> Switches:address
	wire         mm_interconnect_0_sevseg4msb_s1_chipselect;                // mm_interconnect_0:SevSeg4MSB_s1_chipselect -> SevSeg4MSB:chipselect
	wire  [31:0] mm_interconnect_0_sevseg4msb_s1_readdata;                  // SevSeg4MSB:readdata -> mm_interconnect_0:SevSeg4MSB_s1_readdata
	wire   [1:0] mm_interconnect_0_sevseg4msb_s1_address;                   // mm_interconnect_0:SevSeg4MSB_s1_address -> SevSeg4MSB:address
	wire         mm_interconnect_0_sevseg4msb_s1_write;                     // mm_interconnect_0:SevSeg4MSB_s1_write -> SevSeg4MSB:write_n
	wire  [31:0] mm_interconnect_0_sevseg4msb_s1_writedata;                 // mm_interconnect_0:SevSeg4MSB_s1_writedata -> SevSeg4MSB:writedata
	wire         mm_interconnect_0_sdram_s1_chipselect;                     // mm_interconnect_0:SDRAM_s1_chipselect -> SDRAM:az_cs
	wire  [31:0] mm_interconnect_0_sdram_s1_readdata;                       // SDRAM:za_data -> mm_interconnect_0:SDRAM_s1_readdata
	wire         mm_interconnect_0_sdram_s1_waitrequest;                    // SDRAM:za_waitrequest -> mm_interconnect_0:SDRAM_s1_waitrequest
	wire  [24:0] mm_interconnect_0_sdram_s1_address;                        // mm_interconnect_0:SDRAM_s1_address -> SDRAM:az_addr
	wire         mm_interconnect_0_sdram_s1_read;                           // mm_interconnect_0:SDRAM_s1_read -> SDRAM:az_rd_n
	wire   [3:0] mm_interconnect_0_sdram_s1_byteenable;                     // mm_interconnect_0:SDRAM_s1_byteenable -> SDRAM:az_be_n
	wire         mm_interconnect_0_sdram_s1_readdatavalid;                  // SDRAM:za_valid -> mm_interconnect_0:SDRAM_s1_readdatavalid
	wire         mm_interconnect_0_sdram_s1_write;                          // mm_interconnect_0:SDRAM_s1_write -> SDRAM:az_wr_n
	wire  [31:0] mm_interconnect_0_sdram_s1_writedata;                      // mm_interconnect_0:SDRAM_s1_writedata -> SDRAM:az_data
	wire         mm_interconnect_0_keys_s1_chipselect;                      // mm_interconnect_0:KEYS_s1_chipselect -> KEYS:chipselect
	wire  [31:0] mm_interconnect_0_keys_s1_readdata;                        // KEYS:readdata -> mm_interconnect_0:KEYS_s1_readdata
	wire   [1:0] mm_interconnect_0_keys_s1_address;                         // mm_interconnect_0:KEYS_s1_address -> KEYS:address
	wire         mm_interconnect_0_keys_s1_write;                           // mm_interconnect_0:KEYS_s1_write -> KEYS:write_n
	wire  [31:0] mm_interconnect_0_keys_s1_writedata;                       // mm_interconnect_0:KEYS_s1_writedata -> KEYS:writedata
	wire         mm_interconnect_0_timer_0_s1_chipselect;                   // mm_interconnect_0:timer_0_s1_chipselect -> timer_0:chipselect
	wire  [15:0] mm_interconnect_0_timer_0_s1_readdata;                     // timer_0:readdata -> mm_interconnect_0:timer_0_s1_readdata
	wire   [2:0] mm_interconnect_0_timer_0_s1_address;                      // mm_interconnect_0:timer_0_s1_address -> timer_0:address
	wire         mm_interconnect_0_timer_0_s1_write;                        // mm_interconnect_0:timer_0_s1_write -> timer_0:write_n
	wire  [15:0] mm_interconnect_0_timer_0_s1_writedata;                    // mm_interconnect_0:timer_0_s1_writedata -> timer_0:writedata
	wire         mm_interconnect_0_timer_1_s1_chipselect;                   // mm_interconnect_0:timer_1_s1_chipselect -> timer_1:chipselect
	wire  [15:0] mm_interconnect_0_timer_1_s1_readdata;                     // timer_1:readdata -> mm_interconnect_0:timer_1_s1_readdata
	wire   [2:0] mm_interconnect_0_timer_1_s1_address;                      // mm_interconnect_0:timer_1_s1_address -> timer_1:address
	wire         mm_interconnect_0_timer_1_s1_write;                        // mm_interconnect_0:timer_1_s1_write -> timer_1:write_n
	wire  [15:0] mm_interconnect_0_timer_1_s1_writedata;                    // mm_interconnect_0:timer_1_s1_writedata -> timer_1:writedata
	wire         irq_mapper_receiver0_irq;                                  // JTAG_UART:av_irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                  // KEYS:irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver2_irq;                                  // timer_0:irq -> irq_mapper:receiver2_irq
	wire         irq_mapper_receiver3_irq;                                  // timer_1:irq -> irq_mapper:receiver3_irq
	wire  [31:0] processor_d_irq_irq;                                       // irq_mapper:sender_irq -> Processor:d_irq
	wire         rst_controller_reset_out_reset;                            // rst_controller:reset_out -> [GREEN_LEDs:reset_n, JTAG_UART:rst_n, KEYS:reset_n, On_Chip_Mem:reset, Processor:reset_n, RED_LEDs:reset_n, SDRAM:reset_n, SYSID:reset_n, SevSeg4MSB:reset_n, SevSegment_4LSB:reset_n, Switches:reset_n, irq_mapper:reset, mm_interconnect_0:Processor_reset_n_reset_bridge_in_reset_reset, rst_translator:in_reset, timer_0:reset_n, timer_1:reset_n]
	wire         rst_controller_reset_out_reset_req;                        // rst_controller:reset_req -> [On_Chip_Mem:reset_req, Processor:reset_req, rst_translator:reset_req_in]
	wire         processor_jtag_debug_module_reset_reset;                   // Processor:jtag_debug_module_resetrequest -> rst_controller:reset_in0
	wire         clk_reset_source_reset;                                    // CLK:reset_source_reset -> rst_controller:reset_in1

	QsysSystem_CLK clk (
		.ref_clk_clk        (clk_clk),                //      ref_clk.clk
		.ref_reset_reset    (reset_reset),            //    ref_reset.reset
		.sys_clk_clk        (clk_sys_clk_clk),        //      sys_clk.clk
		.sdram_clk_clk      (sdram_clk_clk),          //    sdram_clk.clk
		.reset_source_reset (clk_reset_source_reset)  // reset_source.reset
	);

	QsysSystem_GREEN_LEDs green_leds (
		.clk        (clk_sys_clk_clk),                            //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address    (mm_interconnect_0_green_leds_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_green_leds_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_green_leds_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_green_leds_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_green_leds_s1_readdata),   //                    .readdata
		.out_port   (green_leds_external_connection_export)       // external_connection.export
	);

	QsysSystem_JTAG_UART jtag_uart (
		.clk            (clk_sys_clk_clk),                                           //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                           //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                   //               irq.irq
	);

	QsysSystem_KEYS keys (
		.clk        (clk_sys_clk_clk),                      //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_keys_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_keys_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_keys_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_keys_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_keys_s1_readdata),   //                    .readdata
		.in_port    (keys_external_connection_export),      // external_connection.export
		.irq        (irq_mapper_receiver1_irq)              //                 irq.irq
	);

	QsysSystem_On_Chip_Mem on_chip_mem (
		.clk        (clk_sys_clk_clk),                             //   clk1.clk
		.address    (mm_interconnect_0_on_chip_mem_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_on_chip_mem_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_on_chip_mem_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_on_chip_mem_s1_write),      //       .write
		.readdata   (mm_interconnect_0_on_chip_mem_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_on_chip_mem_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_on_chip_mem_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),              // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),          //       .reset_req
		.freeze     (1'b0)                                         // (terminated)
	);

	QsysSystem_Processor processor (
		.clk                                   (clk_sys_clk_clk),                                           //                       clk.clk
		.reset_n                               (~rst_controller_reset_out_reset),                           //                   reset_n.reset_n
		.reset_req                             (rst_controller_reset_out_reset_req),                        //                          .reset_req
		.d_address                             (processor_data_master_address),                             //               data_master.address
		.d_byteenable                          (processor_data_master_byteenable),                          //                          .byteenable
		.d_read                                (processor_data_master_read),                                //                          .read
		.d_readdata                            (processor_data_master_readdata),                            //                          .readdata
		.d_waitrequest                         (processor_data_master_waitrequest),                         //                          .waitrequest
		.d_write                               (processor_data_master_write),                               //                          .write
		.d_writedata                           (processor_data_master_writedata),                           //                          .writedata
		.d_readdatavalid                       (processor_data_master_readdatavalid),                       //                          .readdatavalid
		.jtag_debug_module_debugaccess_to_roms (processor_data_master_debugaccess),                         //                          .debugaccess
		.i_address                             (processor_instruction_master_address),                      //        instruction_master.address
		.i_read                                (processor_instruction_master_read),                         //                          .read
		.i_readdata                            (processor_instruction_master_readdata),                     //                          .readdata
		.i_waitrequest                         (processor_instruction_master_waitrequest),                  //                          .waitrequest
		.i_readdatavalid                       (processor_instruction_master_readdatavalid),                //                          .readdatavalid
		.d_irq                                 (processor_d_irq_irq),                                       //                     d_irq.irq
		.jtag_debug_module_resetrequest        (processor_jtag_debug_module_reset_reset),                   //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (mm_interconnect_0_processor_jtag_debug_module_address),     //         jtag_debug_module.address
		.jtag_debug_module_byteenable          (mm_interconnect_0_processor_jtag_debug_module_byteenable),  //                          .byteenable
		.jtag_debug_module_debugaccess         (mm_interconnect_0_processor_jtag_debug_module_debugaccess), //                          .debugaccess
		.jtag_debug_module_read                (mm_interconnect_0_processor_jtag_debug_module_read),        //                          .read
		.jtag_debug_module_readdata            (mm_interconnect_0_processor_jtag_debug_module_readdata),    //                          .readdata
		.jtag_debug_module_waitrequest         (mm_interconnect_0_processor_jtag_debug_module_waitrequest), //                          .waitrequest
		.jtag_debug_module_write               (mm_interconnect_0_processor_jtag_debug_module_write),       //                          .write
		.jtag_debug_module_writedata           (mm_interconnect_0_processor_jtag_debug_module_writedata),   //                          .writedata
		.no_ci_readra                          ()                                                           // custom_instruction_master.readra
	);

	QsysSystem_RED_LEDs red_leds (
		.clk        (clk_sys_clk_clk),                          //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address    (mm_interconnect_0_red_leds_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_red_leds_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_red_leds_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_red_leds_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_red_leds_s1_readdata),   //                    .readdata
		.out_port   (red_leds_external_connection_export)       // external_connection.export
	);

	QsysSystem_SDRAM sdram (
		.clk            (clk_sys_clk_clk),                          //   clk.clk
		.reset_n        (~rst_controller_reset_out_reset),          // reset.reset_n
		.az_addr        (mm_interconnect_0_sdram_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_sdram_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_sdram_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_sdram_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_sdram_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_sdram_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_sdram_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_sdram_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_sdram_s1_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_wire_addr),                          //  wire.export
		.zs_ba          (sdram_wire_ba),                            //      .export
		.zs_cas_n       (sdram_wire_cas_n),                         //      .export
		.zs_cke         (sdram_wire_cke),                           //      .export
		.zs_cs_n        (sdram_wire_cs_n),                          //      .export
		.zs_dq          (sdram_wire_dq),                            //      .export
		.zs_dqm         (sdram_wire_dqm),                           //      .export
		.zs_ras_n       (sdram_wire_ras_n),                         //      .export
		.zs_we_n        (sdram_wire_we_n)                           //      .export
	);

	QsysSystem_SYSID sysid (
		.clock    (clk_sys_clk_clk),                                //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_control_slave_address)   //              .address
	);

	QsysSystem_SevSeg4MSB sevseg4msb (
		.clk        (clk_sys_clk_clk),                            //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address    (mm_interconnect_0_sevseg4msb_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_sevseg4msb_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_sevseg4msb_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_sevseg4msb_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_sevseg4msb_s1_readdata),   //                    .readdata
		.out_port   (sevseg4msb_external_connection_export)       // external_connection.export
	);

	QsysSystem_SevSeg4MSB sevsegment_4lsb (
		.clk        (clk_sys_clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                 //               reset.reset_n
		.address    (mm_interconnect_0_sevsegment_4lsb_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_sevsegment_4lsb_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_sevsegment_4lsb_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_sevsegment_4lsb_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_sevsegment_4lsb_s1_readdata),   //                    .readdata
		.out_port   (sevsegment_4lsb_external_connection_export)       // external_connection.export
	);

	QsysSystem_Switches switches (
		.clk      (clk_sys_clk_clk),                        //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address  (mm_interconnect_0_switches_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_switches_s1_readdata), //                    .readdata
		.in_port  (switches_external_connection_export)     // external_connection.export
	);

	QsysSystem_timer_0 timer_0 (
		.clk        (clk_sys_clk_clk),                         //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         // reset.reset_n
		.address    (mm_interconnect_0_timer_0_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_0_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_0_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_0_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_0_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver2_irq)                 //   irq.irq
	);

	QsysSystem_timer_0 timer_1 (
		.clk        (clk_sys_clk_clk),                         //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         // reset.reset_n
		.address    (mm_interconnect_0_timer_1_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_1_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_1_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_1_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_1_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver3_irq)                 //   irq.irq
	);

	QsysSystem_mm_interconnect_0 mm_interconnect_0 (
		.CLK_sys_clk_clk                               (clk_sys_clk_clk),                                           //                             CLK_sys_clk.clk
		.Processor_reset_n_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                            // Processor_reset_n_reset_bridge_in_reset.reset
		.Processor_data_master_address                 (processor_data_master_address),                             //                   Processor_data_master.address
		.Processor_data_master_waitrequest             (processor_data_master_waitrequest),                         //                                        .waitrequest
		.Processor_data_master_byteenable              (processor_data_master_byteenable),                          //                                        .byteenable
		.Processor_data_master_read                    (processor_data_master_read),                                //                                        .read
		.Processor_data_master_readdata                (processor_data_master_readdata),                            //                                        .readdata
		.Processor_data_master_readdatavalid           (processor_data_master_readdatavalid),                       //                                        .readdatavalid
		.Processor_data_master_write                   (processor_data_master_write),                               //                                        .write
		.Processor_data_master_writedata               (processor_data_master_writedata),                           //                                        .writedata
		.Processor_data_master_debugaccess             (processor_data_master_debugaccess),                         //                                        .debugaccess
		.Processor_instruction_master_address          (processor_instruction_master_address),                      //            Processor_instruction_master.address
		.Processor_instruction_master_waitrequest      (processor_instruction_master_waitrequest),                  //                                        .waitrequest
		.Processor_instruction_master_read             (processor_instruction_master_read),                         //                                        .read
		.Processor_instruction_master_readdata         (processor_instruction_master_readdata),                     //                                        .readdata
		.Processor_instruction_master_readdatavalid    (processor_instruction_master_readdatavalid),                //                                        .readdatavalid
		.GREEN_LEDs_s1_address                         (mm_interconnect_0_green_leds_s1_address),                   //                           GREEN_LEDs_s1.address
		.GREEN_LEDs_s1_write                           (mm_interconnect_0_green_leds_s1_write),                     //                                        .write
		.GREEN_LEDs_s1_readdata                        (mm_interconnect_0_green_leds_s1_readdata),                  //                                        .readdata
		.GREEN_LEDs_s1_writedata                       (mm_interconnect_0_green_leds_s1_writedata),                 //                                        .writedata
		.GREEN_LEDs_s1_chipselect                      (mm_interconnect_0_green_leds_s1_chipselect),                //                                        .chipselect
		.JTAG_UART_avalon_jtag_slave_address           (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //             JTAG_UART_avalon_jtag_slave.address
		.JTAG_UART_avalon_jtag_slave_write             (mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),       //                                        .write
		.JTAG_UART_avalon_jtag_slave_read              (mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),        //                                        .read
		.JTAG_UART_avalon_jtag_slave_readdata          (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                                        .readdata
		.JTAG_UART_avalon_jtag_slave_writedata         (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                                        .writedata
		.JTAG_UART_avalon_jtag_slave_waitrequest       (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                                        .waitrequest
		.JTAG_UART_avalon_jtag_slave_chipselect        (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  //                                        .chipselect
		.KEYS_s1_address                               (mm_interconnect_0_keys_s1_address),                         //                                 KEYS_s1.address
		.KEYS_s1_write                                 (mm_interconnect_0_keys_s1_write),                           //                                        .write
		.KEYS_s1_readdata                              (mm_interconnect_0_keys_s1_readdata),                        //                                        .readdata
		.KEYS_s1_writedata                             (mm_interconnect_0_keys_s1_writedata),                       //                                        .writedata
		.KEYS_s1_chipselect                            (mm_interconnect_0_keys_s1_chipselect),                      //                                        .chipselect
		.On_Chip_Mem_s1_address                        (mm_interconnect_0_on_chip_mem_s1_address),                  //                          On_Chip_Mem_s1.address
		.On_Chip_Mem_s1_write                          (mm_interconnect_0_on_chip_mem_s1_write),                    //                                        .write
		.On_Chip_Mem_s1_readdata                       (mm_interconnect_0_on_chip_mem_s1_readdata),                 //                                        .readdata
		.On_Chip_Mem_s1_writedata                      (mm_interconnect_0_on_chip_mem_s1_writedata),                //                                        .writedata
		.On_Chip_Mem_s1_byteenable                     (mm_interconnect_0_on_chip_mem_s1_byteenable),               //                                        .byteenable
		.On_Chip_Mem_s1_chipselect                     (mm_interconnect_0_on_chip_mem_s1_chipselect),               //                                        .chipselect
		.On_Chip_Mem_s1_clken                          (mm_interconnect_0_on_chip_mem_s1_clken),                    //                                        .clken
		.Processor_jtag_debug_module_address           (mm_interconnect_0_processor_jtag_debug_module_address),     //             Processor_jtag_debug_module.address
		.Processor_jtag_debug_module_write             (mm_interconnect_0_processor_jtag_debug_module_write),       //                                        .write
		.Processor_jtag_debug_module_read              (mm_interconnect_0_processor_jtag_debug_module_read),        //                                        .read
		.Processor_jtag_debug_module_readdata          (mm_interconnect_0_processor_jtag_debug_module_readdata),    //                                        .readdata
		.Processor_jtag_debug_module_writedata         (mm_interconnect_0_processor_jtag_debug_module_writedata),   //                                        .writedata
		.Processor_jtag_debug_module_byteenable        (mm_interconnect_0_processor_jtag_debug_module_byteenable),  //                                        .byteenable
		.Processor_jtag_debug_module_waitrequest       (mm_interconnect_0_processor_jtag_debug_module_waitrequest), //                                        .waitrequest
		.Processor_jtag_debug_module_debugaccess       (mm_interconnect_0_processor_jtag_debug_module_debugaccess), //                                        .debugaccess
		.RED_LEDs_s1_address                           (mm_interconnect_0_red_leds_s1_address),                     //                             RED_LEDs_s1.address
		.RED_LEDs_s1_write                             (mm_interconnect_0_red_leds_s1_write),                       //                                        .write
		.RED_LEDs_s1_readdata                          (mm_interconnect_0_red_leds_s1_readdata),                    //                                        .readdata
		.RED_LEDs_s1_writedata                         (mm_interconnect_0_red_leds_s1_writedata),                   //                                        .writedata
		.RED_LEDs_s1_chipselect                        (mm_interconnect_0_red_leds_s1_chipselect),                  //                                        .chipselect
		.SDRAM_s1_address                              (mm_interconnect_0_sdram_s1_address),                        //                                SDRAM_s1.address
		.SDRAM_s1_write                                (mm_interconnect_0_sdram_s1_write),                          //                                        .write
		.SDRAM_s1_read                                 (mm_interconnect_0_sdram_s1_read),                           //                                        .read
		.SDRAM_s1_readdata                             (mm_interconnect_0_sdram_s1_readdata),                       //                                        .readdata
		.SDRAM_s1_writedata                            (mm_interconnect_0_sdram_s1_writedata),                      //                                        .writedata
		.SDRAM_s1_byteenable                           (mm_interconnect_0_sdram_s1_byteenable),                     //                                        .byteenable
		.SDRAM_s1_readdatavalid                        (mm_interconnect_0_sdram_s1_readdatavalid),                  //                                        .readdatavalid
		.SDRAM_s1_waitrequest                          (mm_interconnect_0_sdram_s1_waitrequest),                    //                                        .waitrequest
		.SDRAM_s1_chipselect                           (mm_interconnect_0_sdram_s1_chipselect),                     //                                        .chipselect
		.SevSeg4MSB_s1_address                         (mm_interconnect_0_sevseg4msb_s1_address),                   //                           SevSeg4MSB_s1.address
		.SevSeg4MSB_s1_write                           (mm_interconnect_0_sevseg4msb_s1_write),                     //                                        .write
		.SevSeg4MSB_s1_readdata                        (mm_interconnect_0_sevseg4msb_s1_readdata),                  //                                        .readdata
		.SevSeg4MSB_s1_writedata                       (mm_interconnect_0_sevseg4msb_s1_writedata),                 //                                        .writedata
		.SevSeg4MSB_s1_chipselect                      (mm_interconnect_0_sevseg4msb_s1_chipselect),                //                                        .chipselect
		.SevSegment_4LSB_s1_address                    (mm_interconnect_0_sevsegment_4lsb_s1_address),              //                      SevSegment_4LSB_s1.address
		.SevSegment_4LSB_s1_write                      (mm_interconnect_0_sevsegment_4lsb_s1_write),                //                                        .write
		.SevSegment_4LSB_s1_readdata                   (mm_interconnect_0_sevsegment_4lsb_s1_readdata),             //                                        .readdata
		.SevSegment_4LSB_s1_writedata                  (mm_interconnect_0_sevsegment_4lsb_s1_writedata),            //                                        .writedata
		.SevSegment_4LSB_s1_chipselect                 (mm_interconnect_0_sevsegment_4lsb_s1_chipselect),           //                                        .chipselect
		.Switches_s1_address                           (mm_interconnect_0_switches_s1_address),                     //                             Switches_s1.address
		.Switches_s1_readdata                          (mm_interconnect_0_switches_s1_readdata),                    //                                        .readdata
		.SYSID_control_slave_address                   (mm_interconnect_0_sysid_control_slave_address),             //                     SYSID_control_slave.address
		.SYSID_control_slave_readdata                  (mm_interconnect_0_sysid_control_slave_readdata),            //                                        .readdata
		.timer_0_s1_address                            (mm_interconnect_0_timer_0_s1_address),                      //                              timer_0_s1.address
		.timer_0_s1_write                              (mm_interconnect_0_timer_0_s1_write),                        //                                        .write
		.timer_0_s1_readdata                           (mm_interconnect_0_timer_0_s1_readdata),                     //                                        .readdata
		.timer_0_s1_writedata                          (mm_interconnect_0_timer_0_s1_writedata),                    //                                        .writedata
		.timer_0_s1_chipselect                         (mm_interconnect_0_timer_0_s1_chipselect),                   //                                        .chipselect
		.timer_1_s1_address                            (mm_interconnect_0_timer_1_s1_address),                      //                              timer_1_s1.address
		.timer_1_s1_write                              (mm_interconnect_0_timer_1_s1_write),                        //                                        .write
		.timer_1_s1_readdata                           (mm_interconnect_0_timer_1_s1_readdata),                     //                                        .readdata
		.timer_1_s1_writedata                          (mm_interconnect_0_timer_1_s1_writedata),                    //                                        .writedata
		.timer_1_s1_chipselect                         (mm_interconnect_0_timer_1_s1_chipselect)                    //                                        .chipselect
	);

	QsysSystem_irq_mapper irq_mapper (
		.clk           (clk_sys_clk_clk),                //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),       // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),       // receiver3.irq
		.sender_irq    (processor_d_irq_irq)             //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (processor_jtag_debug_module_reset_reset), // reset_in0.reset
		.reset_in1      (clk_reset_source_reset),                  // reset_in1.reset
		.clk            (clk_sys_clk_clk),                         //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),          // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req),      //          .reset_req
		.reset_req_in0  (1'b0),                                    // (terminated)
		.reset_req_in1  (1'b0),                                    // (terminated)
		.reset_in2      (1'b0),                                    // (terminated)
		.reset_req_in2  (1'b0),                                    // (terminated)
		.reset_in3      (1'b0),                                    // (terminated)
		.reset_req_in3  (1'b0),                                    // (terminated)
		.reset_in4      (1'b0),                                    // (terminated)
		.reset_req_in4  (1'b0),                                    // (terminated)
		.reset_in5      (1'b0),                                    // (terminated)
		.reset_req_in5  (1'b0),                                    // (terminated)
		.reset_in6      (1'b0),                                    // (terminated)
		.reset_req_in6  (1'b0),                                    // (terminated)
		.reset_in7      (1'b0),                                    // (terminated)
		.reset_req_in7  (1'b0),                                    // (terminated)
		.reset_in8      (1'b0),                                    // (terminated)
		.reset_req_in8  (1'b0),                                    // (terminated)
		.reset_in9      (1'b0),                                    // (terminated)
		.reset_req_in9  (1'b0),                                    // (terminated)
		.reset_in10     (1'b0),                                    // (terminated)
		.reset_req_in10 (1'b0),                                    // (terminated)
		.reset_in11     (1'b0),                                    // (terminated)
		.reset_req_in11 (1'b0),                                    // (terminated)
		.reset_in12     (1'b0),                                    // (terminated)
		.reset_req_in12 (1'b0),                                    // (terminated)
		.reset_in13     (1'b0),                                    // (terminated)
		.reset_req_in13 (1'b0),                                    // (terminated)
		.reset_in14     (1'b0),                                    // (terminated)
		.reset_req_in14 (1'b0),                                    // (terminated)
		.reset_in15     (1'b0),                                    // (terminated)
		.reset_req_in15 (1'b0)                                     // (terminated)
	);

endmodule
